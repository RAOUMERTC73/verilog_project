// Code your design here
module and_gate( input in1,
                 input in2,
                 output out
               );
  assign out = a & b;
  
  
endmodule
